BZh91AY&SYb�� �_�Px����������P�WG���jA5�$���z"m24�d���Q��z�S@��P5<��" @  h  	OT����@ɧ���   �0`��`ѐ��&��D@��yO&MM4��S0P=@z��4=C�@IoЄ'�BB$���#��``�"!��� %,Ў��1 �8I��oc��"�8409D��k��J-H����̨|�5Z&#�:):d�ҏ���k��S:���2gQ�D�U�D�.E$ƢŖ��+��Z�k�w����O�-���BZ�;�r�s��p��&��r����\F��ק�L����m���ɵ�ޛ��j�Xȳ��C������Mn}Ո.^�������ε��H�"�o��*l,,ꘖ�r�����]<+-JX�Al�-u(��5��Vl6fGO����"�w6���n�&�5T[�,!Cy;���:d���I��pS�Pӳ���a���-�|�KFʮ�26\� 0��fCE�7U�jf|}��*(�%Ua �0{^��,�ڰ,&���c��bd�6� ��W�C	4E�v	�P�d" �d"��(\D	�e�� �0�^�6���;Ye>���F�R�=�1u~�X\�z����(vՆ���!�X�]0M��wk�j��䪁(�:;���Dd�a�YN��q�& ପ���ow����[Rėش�:��=�qh�T;�b�|H�g���[`آ����8�%�"� �����	l�G���������CA(�u���?�}`��[]Z��ec��E �p�~�&� Pb���@��b�sůҜ�,t2Ώ!�����`]��Nv�7kL�l#Z�P���;s)������ڻ}=�e�HX��G̨�yG ��./PH��6��U��Eۯ#�ƭdV��O����	�,��%k!'�9A�̇M��I��Y�8tu���I��A�� f�m�^�d㱑�1:��P�����	
��e$n4�fUId2W=�D��T�(��(Z��E��Ez��0�J.+��Y��� �H]�H{5�	�f�T:X�Ъ�5��vv��篺4��Q���.l���&V�tj٥JҀۭ; ״/��v�̋�,��X�Ej�f
âqTQ�8	5�a���$�I�]	B�ۑM����h���@���9՜�!Q8;��Vj ĝN�9lsiȾ��%�4��8��df�6�b0j�zV�B�,�
�,kY0[*S_˫�/L�����ʵm�[��5���!�D�_��H�
]� 