BZh91AY&SY�pO� �߀Px����������P��/{08�{�]D��$���y�6��i�i��M�P4��5  h     �D
(��G�A��z�� h =M "�$�H����4�1@		��i=A��4��  =CDʽ���R�)@�$c����	HL�Y=�HB*Ў�EZH)���������)m��I\%� ���0°1$ LC�f3�9��(�s����fk_�W?��٧hH�g�r�Dey��C>Ed��S���+2��T�[pТ�x�7 �@� ���*��*k]�lHL��B_Y�ؓҁs���	��Pճam	�]�y�,��`M2���ecK��p�<�-�9�����`�;�Chmt�C���Voph�\r�
��Q@5�ǽ�WJL58�jX#J��C��p�d2�� U5��"L��E�@�
��F��D>���j���1&�P1�fv��h<ܻd�1tm��h ��x�qp�R�b3Tq���;�b��F��ى���@ @x  ci���}��-�o.��1�%ZR������B�Q�H�%�Uh2OD5$�Cj P�Be�ʉ@��-���A�Z3r��@���JNd�g�)��ys[��U�[�u=u|<ꮲ8j��@�Md`��݇�����k�L�-jy�����n/;�|m2�&B�Y�^~��c��dp�N��U�Y ��ӥ����ƴ�I�ؕ�f�O� @��Z��*�f���O�3���TsNA.&��+��0b�(Hz�����ŷ�I��mwk6��OUc�O6����3OWm�tCLs)��ZP�#��(N)�V�%9�̰:��ĥ�3~�#������Xܘ��Mb��V,�Jf�9v����GWL}��@@0J�a
B]�4q��)ܰ�u�"�
���a�A6&Exk&Uvڹ+}6-FhK
oH_�-&BN<I��[��v+�i�V����ȷ ĶP̹�܃�]K˃Qt�L����� ���d�7�3
 ���.݇$
Ui6N"&���dՓã�albPR�;��"��v�86\�Hzs�!�!F���C��}���p8�j^�Ƞ?!���ti�r��-�������e��LBq���$�3�=�/�gk�������(� ��Aݬ��A�vѪc�Wu�ʦdj�|���J����Pwq�օju�ْE9N訰%���
VȘUӎU�b3����L�+�)���\�iHS��UPK)#U�8v@o�5D#�IR�Y+O��3�7H60X�+���H�
�	� 