BZh91AY&SYסv p_�Px����������`����ʹ ��7��"TBH�S�d5<�e1��=A�����i�	)G�4� � �  ���&L�20�&�db``jD��4���h4L��F�����d h   b EA	���h�Se2zFA� ��G�I@
*V���@e��� +B#�Q�D\@��R�,�i�Z$A�S�	(�ޞ��(����u�W�t��T����%"#{K#;��謸a�=�:�sX�9�S�S�x4�$\��%��V΢(M� �����I�x p���@#�����|��`[�)�j�������w�Ou%k�o�K���$�>m�+=23"����di~������*l���������YF!�+w�|tf'�@�{�Y��Z�2UT��!k��K�Ȯ5baë�)_�.�c���A��Y���LI�E��1{ꁒ�'�,hk��I~T+�W]��916d�B;�L\H��N ������ �P]�Çy�DE�I��͒Y����D(,3V�;uHi��c�s%r��.hIͫ�ᣲ!�D�8��S(am C��-�<�Q}-.&�
(���I�v�A2GV��`Q�V� �p�����Uq��Y�͇����Lp�r��r��s�Uͪtקk{!��,jr�G��滍TXq`���$By�F�qP�=�،Nv�ڝ+W��@,�돽Q��ub^��RK�Cǻ[Pu�oS[�$R�L:S�}z"ȇë%�$Y`ܜ�&�@s2�t�b*�ɖ�2 k<,Ź��p�C�V����O:�gf�m�m^n�(�"d�FX��Q�J*�FB��Ԇ�\���c�6�� �찮G39R����Ǔ3��"�r��%�����O���TQ]uV$!(�?V��Dh`�=�a����\�2�a/���FPx����U]H�ƭ.�UX\�*IC	dX�
Vb���EU1e0�Sj�rd`P2Bұ�����8@��A߲O�}9��2˖�Ux��1|��(���\�ݕ�9Il�ȸ���5Ψ�$#?��o���QQ�Æ3 �&BH�Wa���Y����'gJB����s��&��e�Ȕ�(V0�:�"@�B�6°(��MW	u��"?��F*�R�Y��"��q�¨�-V�ޔ��|� ��Cp`�v�V����Y����4A$"]�fP����Ub��XvN1%y$����]��&a|F'���'i]��9����b�����BS0ۗ����Ú��B��%!��;i"޷�bz9a 5�t8�9��6�bU�ʥ�}e3W�p�/�1 ��HrZ��)�c��p_��)d�(������8����暗��Æ������=R�6��'�"ȋ�A'M�6'i��P��� ~2M���lA�C���Y&�� �UP�*f�%�Y�($����7�;/���e���i�����3j�� �'�-�Ӳ3�";�>�s��B;L�D}vv��#հ2�`���%t��u�,ji8L��nBA���FsA��3$���b�P�i���M�����7�� k����c� ���GS�$(��IE�����r ��Dw�ImοQ��|KT#7{;Z�a���.�p�!�B�