BZh91AY&SY��ў �߀Px����������P~w���Th��&����i�2�SF@h�h�hC@�4�QO� P     "h����
Pi��   � 0&&�	�&L�&	���I ����'����@���Q��E=��J�^���3��
?��l"J��i�l�� =0���NkB�������yrs��N��mxW@6�0B��*	O���KÃ�D��.GT�o�x��=��ӝ�'��㍱݀���V�ć�U�}�l�1T�k���ۼ���&���M�Z���)��<_n��g7n����c��-_j����ZZGImmh�_Ebu�`e�2��YB�6ډ1�"�6oawN�㙧r�Ŗ�[����jb��Rݡ�{[ʻ ��I"�.����c�n2��(�(B�f��%IQ����d���2���%h��T��e}BS�B� ��Y��nb�����&��j]��1�@x�����#`=Ch,U!T,1ff(8�FX��'8�S@MKp� й�W*��+3�"���/6��^Is�*�|�Y�66���LB �g.���fd �>!.8�R�Z�NSՈmH���+qI��,8��)D2�o��� ( ��K"��tu��(E�I�k��W�),�Æ:�.x�?��3�]��P���E�R�	0�&Q ��&�5��/�h�|�D��>\�so��~V��L�O��d(�5q���O������|L���7I@$I$I7��	�>A��������Y��T�n���G��K1uW��"o��:&Ͳ���n]7�0s���B�GR�~[����Z��!ø��/�D��Eipn����Z�b<�[�F,"s.�U|u_�( ��cE��[���.����<5��!hrr�I|��	��R�b(}7r!����AEd]��N�X�}�����QA�m�8���3�O��Z��dL�Ivk��!k����̐��QKfⴘ������A,��f���X��\��5$ON�&�b&�݅���-�@<�N!��m���j6�m��:�PHty��,"V �t��h��XD��q9y������-���X���#Q�q+n
���t{B[e���CF�Vc��L�%�Z��ݤ��&�0����f�{1+��ܖ0��x��f5yN74H�g�v��x�ٹ6��D�d�v�xc�G�n]+���`��QN0���)��f��