BZh91AY&SY_�� �_�Px����������P�6�e�њm-HH�SЧ�M4���CS�Ѧ�i��dhhz���2$�    �@  H�$��?SɣQ4�(�����Si�0L@0	�h�h`ba"��䞚��CM4~���� 1 �z�I/�HP��`H��B��B�e0Б)	�ò_��E���]�������{���+Hn�r\�drop���^���42�i�����j���ۗ
&��Yd�z[f���B��i��� �֢�j�,��N�U�Y��kkV�9R��=�M�0� Ƙ$��=�jM۟�!3�}�ZN�E�%��6�g$C��-#9o���-�k.zƌ`���')��5:D�]����ә���[{�!���I��!�B�T΃ӝ�d�k%�f�oT�mV�`���!���i�0�"UF�&���N~t$(RLΎ��0&¹8zn�Tȧ�K�*�I���j@�XMJS(.�(�W�9�:6��9�.��1��/��y$lm�m��i
�m*����K��r��-UP%i�Υ��*D4���6bU4Xq)6���l�adAa���4+`���A`�[6\ն���+���.�ܵ�?j�
��fO�y���i#~/g�����{~7�aɚJ��q
^Bd��s���Hz�ܖ���1��!2��T�Я�u�8<=�h%$���fnVqu?�w�v*?Uh�%"3����k66��1���m��V�
!yR��ś�r��Ƥ's�ܖ�\`�ԌMm��~N#����&;Z�W�B۬����%T��N�PК�C��� a$(��� ����t��I��<�C�����Y�L\l&�l�ɝ��D�6YӋx����6��xY=��`J7�D�JH�4O�e�">l�Q�(��6ו��Q2��r��jX�_,н!h�32p8tI���[c�LS�q��'l�΅�3�]��o�a.fh��$eE0Z�W��%$�2Q�l�E�dWF�($"�"�Q0K��sqJ�-��R�dK2yHU�K��_������z���1�`���=�D|G`�+��D[�\��G#_^��'E%�3 ״0HVHR<�թu�g}�!r���5�M��41Ń��'���ͣ��{kUd�Q����O9��*s��{����jB�9>�h5�H��lTX�0�B�q$@��0��#V�����_�f���P�X�kHR�*���FU��dt�,��dU*eg��3�"+��w$S�	�Q`